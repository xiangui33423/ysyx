module ysyx_23060096_npc (
    input   [31:0] inst,
    output  [31:0] pc
);



endmodule //ysyx_23060096_NPC