`include "decoder.v"
`include "encoder.v"

module top (
    
);

endmodule //top