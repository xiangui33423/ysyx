module ysyx_23060096_NPC (
    
);

endmodule //ysyx_23060096_NPC