module ysyx_23060096_IDU (
    
);

endmodule //ysyx_23060096_IDU