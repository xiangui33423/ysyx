module ysyx_23060096_IFU (
    
);

endmodule //ysyx_23060096_IFU