module ysyx_23060096_EXU (
    
);

endmodule //ysyx_23060096_EXU