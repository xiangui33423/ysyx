module ysyx_23060096_PCreg (
    input         clk,
    input         rst_n,
    input  [31:0] pc,
    input  []
);

endmodule //ysyx_23060096_PCreg