module main (
    input [7:0] data,
    input       ready,
    input       overflow
);



endmodule //main
