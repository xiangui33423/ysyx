module ysyx_23060096_npc (
    input          clk,
    input          rstn,
    input   [31:0] inst,
    output  [31:0] pc
);

//========IF=======



endmodule //ysyx_23060096_NPC